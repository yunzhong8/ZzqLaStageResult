/*
*作者：zzq
*创建时间：2023-03-31
*email:3486829357@qq.com
*github:yunzhong8
*输入：
*输出：
*模块功能：
*
*/
/*************\
bug:
\*************/
`include "DefineModuleBus.h"
module Preif_IF(
    input  wire  clk      ,
    input  wire  rst_n    ,

    input wire preif_to_if_valid_i,
    input wire if_allowin_i,
    output reg if_valid_o,
    input wire excep_flush_i,
    
    input wire  inst_en_i,
    input  wire [`PcWidth]    pc_i           ,
    output reg inst_en_o,
    output wire  [`PiToIfBusWidth]  to_if_obus
);

/***************************************input variable define(输入变量定义)**************************************/

/***************************************output variable define(输出变量定义)**************************************/
reg  [`PcWidth] pc_o;
/***************************************parameter define(常量定义)**************************************/

/***************************************inner variable define(内部变量定义)**************************************/

/****************************************input decode(输入解码)***************************************/


/****************************************output code(输出解码)***************************************/
assign to_if_obus = pc_o;
/*******************************complete logical function (逻辑功能实现)*******************************/
    always@(posedge clk)begin
        if(rst_n==`RstEnable)begin
            pc_o <= 32'h1bff_fffc;
            inst_en_o<=1'b0;
        end else if(preif_to_if_valid_i&& if_allowin_i)begin
            inst_en_o<=inst_en_i;
            pc_o <= pc_i;
        end else begin
           inst_en_o<=inst_en_o;
            pc_o <= pc_o;
        end
        
    end
     always@(posedge clk)begin
        if(rst_n == `RstEnable || excep_flush_i)begin
            if_valid_o <= 1'b0;
        end else if(if_allowin_i)begin
            if_valid_o <= preif_to_if_valid_i;
        end else begin
             if_valid_o <= if_valid_o;
        end
    end
endmodule
